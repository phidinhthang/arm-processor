library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_textio.all;
use std.textio.all;

package util is
	type imemtype is array (natural range <>) of std_logic_vector;
	type dmemtype is array (natural range <>) of std_logic_vector;
end package util;

package body util is

end package body util;
